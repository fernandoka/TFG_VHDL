----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Fernando Candelario Herrero
-- 
-- Create Date: 14.12.2019 20:22:30
-- Design Name: 
-- Module Name: MyDummyDDR2 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.3
-- Additional Comments:
--					 		
--
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity MyDummyDDR2 is
  Port ( 
        rst_n           :   in  std_logic;
        clk             :   in  std_logic;
		addr			:	in	std_logic_vector(22 downto 0);
		cen             :	in	std_logic; -- low to request a read
        rd              :	in	std_logic; -- One cycle low to request a read
        wr              :	in	std_logic; -- One cycle low to request a read
		ack			    :	out	std_logic; -- One cycle high to notify the reception of a new byte
		data_in         :   in std_logic_vector(15 downto 0);
		data_out		:	out	std_logic_vector(127 downto 0)
  );
-- Attributes for debug
--attribute   dont_touch    :   string;
--attribute   dont_touch  of  MidiRom  :   entity  is  "true";
end MyDummyDDR2;

architecture Behavioral of MyDummyDDR2 is
	constant	MAX_ROWS	:	natural	:= 418;
	
	type romType	is array (0 to MAX_ROWS) of std_logic_vector (127 downto 0);
-- 1=>X"ff00081802040458ff00080700006b72",
-- Papermoon.mid
	constant romRd : romType :=(
0=>X"544de00102000100060000006468544d", 1=>X"ff00081802040458ff00080700006b72", 2=>X"000079b0001cc8060351ff0000fe0259", 3=>X"00005d00005b00400a006407b00000c0", 
4=>X"814046190043478340439000000121ff", 5=>X"43638140430d0045638140450d004663", 6=>X"0d0045638140450d0046638140460d00", 7=>X"40450d0046638140460d004363814043", 
8=>X"638140460d0043638140430d00456381", 9=>X"0043638140430d0045638140450d0046", 10=>X"0d004663815246190043478350436d83", 11=>X"55460d0043638154430d004563815345", 
12=>X"638158430d0045638156450d00466381", 13=>X"004563815a450d0046638159460d0043", 14=>X"450d004663815c460d004363815b430d", 15=>X"51ff6d83004363815e430d004563815d", 
16=>X"000046578a5052005046900020a10703", 17=>X"19005900004d4783505900504d490052", 18=>X"00504a31005700004b0f87505700504b", 19=>X"8a505400504831005600004a0f875056", 
20=>X"50560700547150543183005400004857", 21=>X"56478350565785005471505407005671", 22=>X"578a5052005046190051478350511900", 23=>X"00004d4783505900504d490052000046", 
24=>X"31005700004b0f87505700504b190059", 25=>X"00504831005600004a0f87505600504a", 26=>X"3c2e070351ff490054000048578a5054", 27=>X"8200450f875045190046478350469000", 
28=>X"3d0041738840417d8100416381404121", 29=>X"403719003a4783403a31003a0f87403a", 30=>X"4783403a190039478340391900374783", 31=>X"003e0f87403e31003f0f87403f19003a", 
32=>X"3919003a4783403a19003c4783403c31", 33=>X"88403919003a4783403a190039478340", 34=>X"578a403a7d810037638140373d003973", 35=>X"003a6381403a0d003a6381403a49003a", 
36=>X"3f19003e4783403e0d003c6381403c0d", 37=>X"83403e25003f2b85403f0d003f638140", 38=>X"47834041218200390f87403919003e47", 39=>X"31004100003a0f87404100403a190041", 
40=>X"403a31003a0f87403a0d003a6381403a", 41=>X"478340391900374783403719003a4783", 42=>X"85403f00403c19003a4783403a190039", 43=>X"403e0d003e6381403e25003f00003c2b", 
44=>X"4783403a19003c4783403c31003e0f87", 45=>X"003a4783403a1900394783403919003a", 46=>X"3a190037478340373d00397388403919", 47=>X"417d810041638140412d82003a738840", 
48=>X"83403e19003f4783403f190041478340", 49=>X"3e4783403e19003f4783403f19003e47", 50=>X"4783403f00403c19003c4783403c1900", 51=>X"00003a4783403e00403a19003f00003c", 
52=>X"82003e00003a7388403e00403a19003e", 53=>X"3e7d81004100003e6381404100403e2d", 54=>X"3f00403c19004100003e478340410040", 55=>X"4783403e00403a19003f00003c478340", 
56=>X"00003c4783403f00403c19003e00003a", 57=>X"49003e00003a578a403e00403a19003f", 58=>X"432d82003e7388403e19003a4783403a", 59=>X"45005041190046000043478350460050", 
60=>X"82504300503f2d820045000041738850", 61=>X"43578a50460050430b81004300003f55", 62=>X"46000043638150460050434900460000", 63=>X"820045000041738850450050417d8100", 
64=>X"5046190045000041478350450050412d", 65=>X"4500503e3100450f8750453d00467388", 66=>X"6381504600503e19004500003e478350", 67=>X"00003e4783504500503e0d004600003e", 
68=>X"81004600003e6381504600503e190045", 69=>X"5043190048000045478350480050457d", 70=>X"50450050411900460000434783504600", 71=>X"3f4783504300503f1900450000414783", 
72=>X"4100003e7388504100503e1900430000", 73=>X"81004100003e6381504100503e2d8200", 74=>X"503e19004300003f4783504300503f7d", 75=>X"503f00503c19004100003e4783504100", 
76=>X"3e4783504100503e19003f00003c4783", 77=>X"3e00003a7388503e00503a1900410000", 78=>X"81003e00003a6381503e00503a2d8200", 79=>X"503f19003f00003c4783503f00503c7d", 
80=>X"504100503e19004300003f4783504300", 81=>X"3c4783503f00503c19004100003e4783", 82=>X"3e00003a7388503e00503a19003f0000", 83=>X"81003e00003a6381503e00503a2d8200", 
84=>X"3a1582003f00003c2b85503f00503c7d", 85=>X"3c00503925003e00003a2b85503e0050", 86=>X"4783504500503e19003c000039478350", 87=>X"00003e6381504600503e19004500003e", 
88=>X"19004500003e4783504500503e0d0046", 89=>X"50457d81004600003e6381504600503e", 90=>X"50460050431900480000454783504800", 91=>X"41478350450050411900460000434783", 
92=>X"4300003f4783504300503f1900450000", 93=>X"2d82004100003e7388504100503e1900", 94=>X"50417d81004600004363815046005043", 95=>X"450050412d8200450000417388504500", 
96=>X"00450f8750456d830045000041638150", 97=>X"0046738850467d810043638150432182", 98=>X"8350480050467d810046638150462d82", 99=>X"50451900464783504619004800004647", 
100=>X"03905043190046478350461900454783", 101=>X"19004300003f4783504300503f6d0043", 102=>X"00503f0d004600004363815046005043", 103=>X"504100503e7d81004300003f63815043", 
104=>X"4783503f00503c7d81004100003e6381", 105=>X"503a7d81003e6381503e19003f00003c", 106=>X"503e7d81003c6381503c7d81003a6381", 107=>X"638140422d82004200003e7388504200", 
108=>X"0042638140420d0042638140420d0042", 109=>X"3e31003f0f87403f3100410f8740410d", 110=>X"0f87403a61004100003e1f8e40410040", 111=>X"003f1f8e403f31003c0f87403c31003a", 
112=>X"403e00403a00403761003e1f8e403e61", 113=>X"544d002fff01003e00003a0000373f9c", 114=>X"0121ff0000fe0259ff005c0b00006b72", 115=>X"2b0d002b6381502b901e9a7f40b00200", 
116=>X"837f40010040b001502b0d002b638150", 117=>X"6381532d0d002e6381522e19002b9045", 118=>X"002e6381552e0d002b6381542b0d002d", 119=>X"2e0d002b6381582b0d002d6381562d0d", 
120=>X"815b2b0d002d63815a2d0d002e638159", 121=>X"2d63815d2d0d002e63815c2e0d002b63", 122=>X"00502e00502b6d83002b63815e2b0d00", 123=>X"2b903d9c7f40010040b0015037005032", 
124=>X"330050304181003700003200002e0000", 125=>X"3d9c7f40010040b001503c0050360050", 126=>X"502e4181003c00003600003300003090", 127=>X"7f40010040b001503a00503500503200", 
128=>X"4181003a00003500003200002e903d9c", 129=>X"010040b001503500503000502d005029", 130=>X"003500003000002d000029903d9c7f40", 131=>X"40b001403700403200402e00402b4181", 
132=>X"00003200002e00002b903d9c7f400100", 133=>X"01403c00403600403300403041810037", 134=>X"36000033000030903d9c7f40010040b0", 135=>X"3300402e00402b0040274181003c0000", 
136=>X"002b000027903d9c7f40010040b00140", 137=>X"403500403200402e4181003300002e00", 138=>X"00002e901d8e7f40010040b001403a00", 139=>X"3000402d00402961003a000035000032", 
140=>X"0029901d8e7f40010040b00140350040", 141=>X"00403200402b61003500003000002d00", 142=>X"3200002b9045837f40010040b0014037", 143=>X"2b4783403700403200402b1900370000", 
144=>X"403700403200402b1900370000320000", 145=>X"403200402b19003700003200002b4783", 146=>X"402b19003700003200002b4783403700", 147=>X"003700003200002b4783403700403200", 
148=>X"003200002b4783403700403200402b19", 149=>X"002b4783403700403200402b19003700", 150=>X"83403700403200402b19003700003200", 151=>X"00403300403019003700003200002b47", 
152=>X"330000309045837f40010040b0014036", 153=>X"30478340360040330040301900360000", 154=>X"40360040330040301900360000330000", 155=>X"40330040301900360000330000304783", 
156=>X"40301900360000330000304783403600", 157=>X"00360000330000304783403600403300", 158=>X"00330000304783403600403300403019", 159=>X"00304783403600403300403019003600", 
160=>X"83403600403300403019003600003300", 161=>X"00402e00402719003600003300003047", 162=>X"2e0000279045837f40010040b0014033", 163=>X"274783403300402e0040271900330000", 
164=>X"403300402e00402719003300002e0000", 165=>X"402e00402719003300002e0000274783", 166=>X"402719003300002e0000274783403300", 167=>X"003300002e0000274783403300402e00", 
168=>X"002e0000274783403300402e00402719", 169=>X"00274783403300402e00402719003300", 170=>X"83403300402e00402719003300002e00", 171=>X"00403000402919003300002e00002747", 
172=>X"300000299045837f40010040b0014035", 173=>X"29478340350040300040291900350000", 174=>X"40350040300040291900350000300000", 175=>X"40300040291900350000300000294783", 
176=>X"40291900350000300000294783403500", 177=>X"00350000300000294783403500403000", 178=>X"00300000294783403500403000402919", 179=>X"00294783403500403000402919003500", 
180=>X"83403500403000402919003500003000", 181=>X"00402e00402719003500003000002947", 182=>X"2e0000279045837f40010040b0014033", 183=>X"274783403300402e0040271900330000", 
184=>X"403300402e00402719003300002e0000", 185=>X"402e00402719003300002e0000274783", 186=>X"402919003300002e0000274783403300", 187=>X"9045837f40010040b001403500403000", 
188=>X"35004030004029190035000030000029", 189=>X"30004029190035000030000029478340", 190=>X"29190035000030000029478340350040", 191=>X"35000030000029478340350040300040", 
192=>X"40010040b001403700403200402b1900", 193=>X"00402b19003700003200002b9045837f", 194=>X"19003700003200002b47834037004032", 195=>X"00003200002b4783403700403200402b", 
196=>X"00002b4783403700403200402b190037", 197=>X"4783403700403200402b190037000032", 198=>X"3700403200402b19003700003200002b", 199=>X"3200402b19003700003200002b478340", 
200=>X"2b19003700003200002b478340370040", 201=>X"3700003200002b478350370050320050", 202=>X"40010040b001503300502e0050271900", 203=>X"00502719003300002e0000279045837f", 
204=>X"19003300002e0000274783503300502e", 205=>X"00002e0000274783503300502e005027", 206=>X"0000274783503300502e005027190033", 207=>X"4783503300502e00502719003300002e", 
208=>X"3300502e00502719003300002e000027", 209=>X"2e00502719003300002e000027478350", 210=>X"2719003300002e000027478350330050", 211=>X"3300002e0000274783503300502e0050", 
212=>X"40010040b00150350050300050291900", 213=>X"0050291900350000300000299045837f", 214=>X"19003500003000002947835035005030", 215=>X"00003000002947835035005030005029", 
216=>X"00002947835035005030005029190035", 217=>X"1f8e5035005030005029190035000030", 218=>X"3700503200502b610035000030000029", 219=>X"003200002b9029857f40010040b00150", 
220=>X"002b2b85503700503200502b25003700", 221=>X"83503700503200502b25003700003200", 222=>X"00502e00502719003700003200002b47", 223=>X"2e0000279029857f40010040b0015033", 
224=>X"272b85503300502e0050272500330000", 225=>X"503300502e00502725003300002e0000", 226=>X"503500502e19003300002e0000274783", 227=>X"00002e9029857f40010040b001503a00", 
228=>X"2b85503a00503500502e25003a000035", 229=>X"3a00503500502e25003a00003500002e", 230=>X"3000502919003a00003500002e478350", 231=>X"00299029857f40010040b00150350050", 
232=>X"85503500503000502925003500003000", 233=>X"0050300050292500350000300000292b", 234=>X"00502b19003500003000002947835035", 235=>X"2b9029857f40010040b0015037005032", 
236=>X"503700503200502b2500370000320000", 237=>X"503200502b25003700003200002b2b85", 238=>X"502719003700003200002b4783503700", 239=>X"9029857f40010040b001503300502e00", 
240=>X"3300502e00502725003300002e000027", 241=>X"2e00502725003300002e0000272b8550", 242=>X"2e19003300002e000027478350330050", 243=>X"29857f40010040b001503a0050350050", 
244=>X"00503500502e25003a00003500002e90", 245=>X"00502e25003a00003500002e2b85503a", 246=>X"19003a00003500002e4783503a005035", 247=>X"857f40010040b0015035005030005029", 
248=>X"50300050292500350000300000299029", 249=>X"50292500350000300000292b85503500", 250=>X"00350000300000294783503500503000", 251=>X"7f40010040b001503700503200502b19", 
252=>X"3200502b25003700003200002b902985", 253=>X"2b25003700003200002b2b8550370050", 254=>X"3700003200002b478350370050320050", 255=>X"40010040b001503300502e0050271900", 
256=>X"00502725003300002e0000279029857f", 257=>X"25003300002e0000272b85503300502e", 258=>X"00002e0000274783503300502e005027", 259=>X"010040b001503a00503500502e190033", 
260=>X"502e25003a00003500002e9029857f40", 261=>X"003a00003500002e2b85503a00503500", 262=>X"003500002e4783503a00503500502e25", 263=>X"0040b001503500503000502919003a00", 
264=>X"292500350000300000299029857f4001", 265=>X"350000300000292b8550350050300050", 266=>X"30000029478350350050300050292500", 267=>X"40b001503700503200502b1900350000", 
268=>X"25003700003200002b9029857f400100", 269=>X"00003200002b2b85503700503200502b", 270=>X"00002b4783503700503200502b250037", 271=>X"b001503300502e005027190037000032", 
272=>X"003300002e0000279029857f40010040", 273=>X"002e0000272b85503300502e00502725", 274=>X"00274783503300502e00502725003300", 275=>X"01503c00503300503019003300002e00", 
276=>X"3c000033000030903d9c7f40010040b0", 277=>X"010040b001503300502e005027418100", 278=>X"502719003300002e0000279045837f40", 279=>X"003300002e0000274783503300502e00", 
280=>X"002e0000274783503300502e00502719", 281=>X"00274783503300502e00502719003300", 282=>X"83503300502e00502719003300002e00", 283=>X"00502e00502719003300002e00002747", 
284=>X"00502719003300002e00002747835033", 285=>X"19003300002e0000274783503300502e", 286=>X"00002e0000274783503300502e005027", 287=>X"b001503c005036005033005030190033", 
288=>X"0036000033000030903d9c7f40010040", 289=>X"403700403200402e00402b4181003c00", 290=>X"00002e00002b903d9c7f40010040b001", 291=>X"00403600403300403041810037000032", 
292=>X"33000030903d9c7f40010040b001403c", 293=>X"2600402200401f4181003c0000360000", 294=>X"001f903d9c7f40010040b001402b0040", 295=>X"ff010040b04181002b00002600002200", 
296=>X"ff010040b04181002b0000260000002f",-- End of Papermoon.mid

297=>X"f4ffeefff4fff1fff4fff5fff4fff9ff",-- 8Sound samples
298=>X"2b00300039003e004100490049005000",

-- OneDividedByDivision Constants
299=>X"00040000000555550008000000100000", 
300=>X"00020000000249250002aaab00033333", 301=>X"000155550001745d0001999a0001c71c", 302=>X"00010000000111110001249200013b14", 303=>X"0000cccd0000d7940000e38e0000f0f1", 304=>X"0000aaab0000b2160000ba2f0000c30c", 
305=>X"00009249000097b400009d8a0000a3d7", 306=>X"00008000000084210000888900008d3e", 307=>X"000071c7000075070000787800007c1f", 308=>X"000066660000690700006bca00006eb4", 309=>X"00005d1700005f4100006186000063e7", 
310=>X"00005555000057260000590b00005b06", 311=>X"00004ec500005050000051ec00005398", 312=>X"0000492500004a7900004bda00004d48", 313=>X"000044440000456c0000469f000047dc", 314=>X"00004000000041040000421100004326", 
315=>X"00003c3c00003d2200003e1000003f04", 316=>X"000038e4000039b100003a8400003b5d", 317=>X"000035e50000369d0000375a0000381c", 318=>X"00003333000033d90000348300003532", 319=>X"000030c300003159000031f400003291", 
320=>X"00002e8c00002f1500002fa100003030", 321=>X"00002c8600002d0300002d8300002e06", 322=>X"00002aab00002b1e00002b9300002c0b", 323=>X"000028f600002960000029cc00002a3a", 324=>X"00002762000027c4000028280000288e", 
325=>X"000025ed00002648000026a400002702", 326=>X"00002492000024e70000253d00002594", 327=>X"0000234f0000239e000023ee0000243f", 328=>X"000022220000226c000022b600002302", 329=>X"000021080000214d00002193000021da", 
330=>X"000020000000204100002082000020c5", 331=>X"00001f0800001f4400001f8200001fc0", 332=>X"00001e1e00001e5700001e9100001ecc", 333=>X"00001d4200001d7800001dae00001de6", 334=>X"00001c7200001ca500001cd800001d0d", 
335=>X"00001bad00001bdd00001c0e00001c40", 336=>X"00001af300001b2000001b4f00001b7d", 337=>X"00001a4200001a6d00001a9900001ac5", 338=>X"0000199a000019c3000019ed00001a17", 339=>X"000018fa000019210000194900001971", 
340=>X"0000186200001887000018ad000018d3", 341=>X"000017d0000017f4000018180000183d", 342=>X"00001746000017680000178a000017ad", 343=>X"000016c1000016e20000170300001724", 344=>X"000016430000166200001681000016a1", 
345=>X"000015ca000015e70000160600001624", 346=>X"00001555000015720000158f000015ac", 347=>X"000014e6000015010000151d00001539", 348=>X"0000147b00001495000014b0000014cb", 349=>X"000014140000142d0000144700001461", 
350=>X"000013b1000013ca000013e2000013fb", 351=>X"000013520000136a0000138100001399", 352=>X"000012f70000130d000013240000133b", 353=>X"0000129e000012b4000012ca000012e0", 354=>X"000012490000125e0000127300001289", 
355=>X"000011f70000120b0000122000001234", 356=>X"000011a8000011bb000011cf000011e3", 357=>X"0000115b0000116e0000118100001194", 358=>X"00001111000011230000113600001148", 359=>X"000010c9000010db000010ed000010ff", 
360=>X"0000108400001095000010a7000010b8", 361=>X"00001041000010520000106200001073", 362=>X"00001000000010100000102000001031", 363=>X"00000fc100000fd100000fe000000ff0", 364=>X"00000f8400000f9300000fa200000fb2", 
365=>X"00000f4900000f5700000f6600000f75", 366=>X"00000f0f00000f1d00000f2c00000f3a", 367=>X"00000ed700000ee500000ef300000f01", 368=>X"00000ea100000eae00000ebc00000ec9", 369=>X"00000e6c00000e7900000e8600000e94", 
370=>X"00000e3900000e4600000e5200000e5f", 371=>X"00000e0700000e1300000e2000000e2c", 372=>X"00000dd600000de200000def00000dfb", 373=>X"00000da700000db300000dbf00000dcb", 374=>X"00000d7900000d8500000d9000000d9c", 
375=>X"00000d4c00000d5800000d6300000d6e", 376=>X"00000d2100000d2c00000d3700000d41", 377=>X"00000cf600000d0100000d0b00000d16", 378=>X"00000ccd00000cd700000ce100000cec", 379=>X"00000ca400000cae00000cb800000cc3", 
380=>X"00000c7d00000c8700000c9000000c9a", 381=>X"00000c5600000c6000000c6a00000c73", 382=>X"00000c3100000c3a00000c4300000c4d", 383=>X"00000c0c00000c1500000c1e00000c28", 384=>X"00000be800000bf100000bfa00000c03", 
385=>X"00000bc500000bce00000bd700000bdf", 386=>X"00000ba300000bab00000bb400000bbd", 387=>X"00000b8100000b8a00000b9200000b9a", 388=>X"00000b6100000b6900000b7100000b79", 389=>X"00000b4100000b4900000b5100000b59", 
390=>X"00000b2100000b2900000b3100000b39", 391=>X"00000b0300000b0a00000b1200000b1a", 392=>X"00000ae500000aec00000af400000afb", 393=>X"00000ac700000acf00000ad600000add", 394=>X"00000aab00000ab200000ab900000ac0", 
395=>X"00000a8f00000a9500000a9d00000aa4", 396=>X"00000a7300000a7a00000a8100000a88", 397=>X"00000a5800000a5f00000a6500000a6c", 398=>X"00000a3d00000a4400000a4b00000a51", 399=>X"00000a2300000a2a00000a3000000a37", 
400=>X"00000a0a00000a1000000a1700000a1d", 401=>X"000009f1000009f7000009fe00000a04", 402=>X"000009d9000009df000009e5000009eb", 403=>X"000009c1000009c7000009cd000009d3", 404=>X"000009a9000009af000009b5000009bb", 
405=>X"00000992000009980000099d000009a3", 406=>X"0000097b00000981000009870000098c", 407=>X"000009650000096b0000097000000976", 408=>X"0000094f000009550000095a0000095f", 409=>X"0000093a0000093f000009440000094a", 
410=>X"000009250000092a0000092f00000934", 411=>X"00000910000009150000091a0000091f", 412=>X"000008fc00000901000009060000090b", 413=>X"000008e8000008ec000008f1000008f6", 414=>X"000008d4000008d9000008de000008e3", 
415=>X"000008c1000008c5000008ca000008cf", 416=>X"000008ae000008b2000008b7000008bc", 417=>X"0000089b000008a0000008a4000008a9", 418=>X"000008890000088d0000089200000896"
);

begin

process(rst_n,clk,rd,wr,addr)
	variable regVal	:	std_logic_vector(127 downto 0);
	variable romWr : std_logic_vector (15 downto 0);	
begin
    
	data_out <= regVal;
	
    if rst_n='0' then
		regVal :=(others=>'0');
		ack <='0';
		
    elsif rising_edge(clk) then
		ack <='0';
		if cen='0' and (wr='0' or rd='0') then
            ack <='1'; --
            if unsigned(addr) < MAX_ROWS then
                if wr='0' then
                    romWr := data_in;
                elsif rd='0' then
                    regVal := romRd(to_integer(unsigned(addr)));
                end if;
            end if;
            
       end if;--cen='0'		
	end if;
end process;
  
end Behavioral;
